`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:58:36 08/17/2014 
// Design Name: 
// Module Name:    PUF_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PUF_unit #(parameter N_CB = 64, N = 16)(
    input wire in,
	 input wire [N_CB-1:0] challenge,
	 input wire [N-1:0] tune,
    output wire out
    );


endmodule
